`timescale 1ns/1ps

`include "Rx.v"

module TB();

  reg clk;
  reg enb;
  reg reset;
  reg L0;
  reg L1;
  reg L2;
  reg L3;

  wire [3:0] S;
  wire [7:0] data;

  Rx prueba(.clk(clk), .enb(enb), .reset(reset), .L0(L0), .L1(L1), .L2(L2), .L3(L3), .S(S), .data(data));

  always #1 clk = !clk;

  initial begin
  $display ("test");
  $dumpfile("gtkws/testRx.vcd");
  $dumpvars;
  $display ("time\t    clk  , data  ,   enb  ,   S   ,   L0  ,   L1  ,   L2  ,   L3 ");
  $monitor ("%g\t      %b     %h       %b      %b        %b       %b       %b      %b",
  $time, clk, data, enb, S, L0, L1, L2, L3);

  clk <= 0;
  reset <= 1'b1;
  enb <= 0;
  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;

  # 4
  @ (posedge clk);
  reset <= 1'b0;
  enb <= 1;


  # 4
      $display("inicio");


  // IDLE
  @ (posedge clk);
  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

//COM

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  //STP

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 0;
  L1 <= 1;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  //DATA=00000001
  L0 <= 1;
  L1 <= 0;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 0;
  L3 <= 0;
  # 1

  //DATA=00000010
  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 1;
  L3 <= 0;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 0;
  L3 <= 0;
  # 1

  //END
  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 0;
  L1 <= 0;
  L2 <= 0;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 0;
  L2 <= 1;
  L3 <= 1;
  # 1

  L0 <= 1;
  L1 <= 1;
  L2 <= 0;
  L3 <= 1;
  # 64







  $finish;
  end



endmodule
